LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; --use CONV_INTEGER

ENTITY fetch IS
 PORT  (
  PC: IN STD_LOGIC_VECTOR(31 downto 0);  -- Program Counter
  Instruction: OUT STD_LOGIC_VECTOR(31 downto 0)   -- Instruction
  );
END fetch;

ARCHITECTURE rtl OF fetch IS
  
  TYPE rom IS ARRAY (0 TO 1339) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
  
  -- Instruction Memory
  -- Big Endian
  CONSTANT imem: 
  rom:=rom'(
				
				
--				"00000100", "00000011", "11101110", "11011011", --32--addi
--				"00010100", "01100011", "00000000", "00010000", --36--shl
--				"00000100", "00000101", "10100101", "00100001", --32--addi 
--				"00010100", "10100101", "00000000", "00010000", --36--shl
--				"00011000", "10100101", "00000000", "00010000", --36--shr
--				"00000000", "01100101", "00011000", "00010011", --40--or
--				"00100000", "00000011", "00000000", "00101110", --44d0--eedba521--56
				
--				"00000100", "00000011", "11101110", "11011011", --32--addi
--				"00010100", "01100011", "00000000", "00010000", --36--shl
--				"00000100", "00000101", "10100101", "00100001", --32--addi r0 r5 0xa521
--				"00010100", "10100101", "00000000", "00010000", --36--shl
--				"00011000", "10100101", "00000000", "00010000", --36--shr
--				"00000000", "01100101", "00011000", "00010011", --40--or
				
				"11111100", "00000000", "00000000", "00000000", --  addr 0 Halt
				"11111100", "00000000", "00000000", "00000000",
				
				"00000000", "00000000", "00000000", "00000000", --08 
			   "00000000", "00000000", "00000000", "00000000",	--12
				"00000000", "00000000", "00000000", "00000000",	--16
				"00000000", "00000000", "00000000", "00000000", --20	
				"00000000", "00000000", "00000000", "00000000",	--24
				"00000000", "00000000", "00000000", "00000000", --28
				"00000000", "00000000", "00000000", "00000000",	--32
				"00000000", "00000000", "00000000", "00000000", --36
				
				
				"00000000", "00000000", "00000000", "00000000",	--40
				"00000000", "00000000", "00000000", "00000000",	--44
				"00000000", "00000000", "00000000", "00000000",	--48
				"00000000", "00000000", "00000000", "00000000",	--52
				"00000000", "00000000", "00000000", "00000000",	--56
				"00000000", "00000000", "00000000", "00000000",	--60
				"00000000", "00000000", "00000000", "00000000",	--64
				"00000000", "00000000", "00000000", "00000000",	--68
				"00000000", "00000000", "00000000", "00000000",	--72
				"00000000", "00000000", "00000000", "00000000", --76	
				
				
				"00000000", "00000000", "00000000", "00000000",	--80
				"00000000", "00000000", "00000000", "00000000",	--84
				"00000000", "00000000", "00000000", "00000000",	--88
				"00000000", "00000000", "00000000", "00000000",	--92
				"00000000", "00000000", "00000000", "00000000",	--96
				"00000000", "00000000", "00000000", "00000000",	--100
				"00000000", "00000000", "00000000", "00000000", --104	
				
				"00000000", "00000000", "00000000", "00000000",	--108
				"00000000", "00000000", "00000000", "00000000",	--112
				"00000000", "00000000", "00000000", "00000000",	--116
				"00000000", "00000000", "00000000", "00000000",	--120
				"00000000", "00000000", "00000000", "00000000",	--124
				"00000000", "00000000", "00000000", "00000000",	--128
				"00000000", "00000000", "00000000", "00000000",	--132
				"00000000", "00000000", "00000000", "00000000",	--136
				"00000000", "00000000", "00000000", "00000000",	--140
				"00000000", "00000000", "00000000", "00000000", -- 144	
				
				"00000000", "00000000", "00000000", "00000000",	--148
				"00000000", "00000000", "00000000", "00000000",	--152
				"00000000", "00000000", "00000000", "00000000",	--156
				"00000000", "00000000", "00000000", "00000000",	--160
				"00000000", "00000000", "00000000", "00000000",	--164
				"00000000", "00000000", "00000000", "00000000",	--168
				"00000000", "00000000", "00000000", "00000000",	--172
				"00000000", "00000000", "00000000", "00000000",	--176
				"00000000", "00000000", "00000000", "00000000",	--180
				"00000000", "00000000", "00000000", "00000000", -- 184	
				
				"00000000", "00000000", "00000000", "00000000",	--188
				"00000000", "00000000", "00000000", "00000000",	--192
				"00000000", "00000000", "00000000", "00000000",	--196
				"00000000", "00000000", "00000000", "00000000",	--200
				"00000000", "00000000", "00000000", "00000000",	--204
				"00000000", "00000000", "00000000", "00000000",	--208
				"00000000", "00000000", "00000000", "00000000",	--212
				"00000000", "00000000", "00000000", "00000000",	--216
				"00000000", "00000000", "00000000", "00000000",	--220
				"00000000", "00000000", "00000000", "00000000", --224	
				
				"00000000", "00000000", "00000000", "00000000",	--228
				"00000000", "00000000", "00000000", "00000000",	--232
				"00000000", "00000000", "00000000", "00000000",	--236
				"00000000", "00000000", "00000000", "00000000",	--240
				"00000000", "00000000", "00000000", "00000000",	--244
				"00000000", "00000000", "00000000", "00000000",	--248
				"00000000", "00000000", "00000000", "00000000",	--252
				"00000000", "00000000", "00000000", "00000000",	--256
				"00000000", "00000000", "00000000", "00000000",	--260
				"00000000", "00000000", "00000000", "00000000", --264 
				
				"00000000", "00000000", "00000000", "00000000",	--268
				"00000000", "00000000", "00000000", "00000000",	--272
				"00000000", "00000000", "00000000", "00000000",	--276
				"00000000", "00000000", "00000000", "00000000",	--280
				"00000000", "00000000", "00000000", "00000000",	--284
				"00000000", "00000000", "00000000", "00000000",	--288
				"00000000", "00000000", "00000000", "00000000",	--292
				"00000000", "00000000", "00000000", "00000000",	--296
				"00000000", "00000000", "00000000", "00000000",	--300
				"00000000", "00000000", "00000000", "00000000", --304 
				
				"00000000", "00000000", "00000000", "00000000",	--308
				"00000000", "00000000", "00000000", "00000000",	--312
				"00000000", "00000000", "00000000", "00000000",	--316
				"00000000", "00000000", "00000000", "00000000",	--320
				"00000000", "00000000", "00000000", "00000000",	--324
				"00000000", "00000000", "00000000", "00000000",	--328
				"00000000", "00000000", "00000000", "00000000",	--332
				"00000000", "00000000", "00000000", "00000000",	--336
				"00000000", "00000000", "00000000", "00000000",	--340
				"00000000", "00000000", "00000000", "00000000", --344	
				
				"00000000", "00000000", "00000000", "00000000",	--348
				"00000000", "00000000", "00000000", "00000000",	--352
				"00000000", "00000000", "00000000", "00000000",	--356
				"00000000", "00000000", "00000000", "00000000",	--360
				"00000000", "00000000", "00000000", "00000000",	--364
				"00000000", "00000000", "00000000", "00000000",	--368
				"00000000", "00000000", "00000000", "00000000",	--372
				"00000000", "00000000", "00000000", "00000000",	--376
				"00000000", "00000000", "00000000", "00000000",	--380
				"00000000", "00000000", "00000000", "00000000", --384 
				
				"00000000", "00000000", "00000000", "00000000",	--388
				"00000000", "00000000", "00000000", "00000000",	--392
				"00000000", "00000000", "00000000", "00000000",	--396
				"00000000", "00000000", "00000000", "00000000",	--400
				"00000000", "00000000", "00000000", "00000000",	--404
				"00000000", "00000000", "00000000", "00000000",	--408
				"00000000", "00000000", "00000000", "00000000",	--412
				"00000000", "00000000", "00000000", "00000000",	--416
				"00000000", "00000000", "00000000", "00000000",	--420
				"00000000", "00000000", "00000000", "00000000", --424 
				
				"00000000", "00000000", "00000000", "00000000",	--428
				"00000000", "00000000", "00000000", "00000000",	--432
				"00000000", "00000000", "00000000", "00000000",	--436
				"00000000", "00000000", "00000000", "00000000",	--440
				"00000000", "00000000", "00000000", "00000000",	--444
				"00000000", "00000000", "00000000", "00000000",	--448
				"00000000", "00000000", "00000000", "00000000",	--452
				"00000000", "00000000", "00000000", "00000000",	--456
				"00000000", "00000000", "00000000", "00000000",	--460
				"00000000", "00000000", "00000000", "00000000", --464 
				
			
				
																				-- Keygen begins
				"00000100", "00000001", "10110111", "11100001", --468
				"00010100", "00100001", "00000000", "00010000", --472
				"00010000", "00100001", "01010001", "01100011", --476
				"00100000", "00000001", "00000000", "00001110", --480
				"00000100", "00000010", "10011110", "00110111", --484
				"00010100", "01000010", "00000000", "00010000", --488
				"00010000", "01000010", "01111001", "10111001", --492
				"00100000", "00000010", "00000000", "00001111", --496
																				-- Keygen begins
				"00011100", "00000001", "00000000", "00001110", --500 
				"00011100", "00000010", "00000000", "00001111", --504
				"00000100", "00000100", "00000000", "00010100", --508
				"00100000", "10000001", "00000000", "00000000", --512
				"00000100", "00000110", "00000000", "00011001", --516
				"00000000", "10000110", "00111000", "00010000", --520
				"00000100", "10000100", "00000000", "00000001", --524
				"00011100", "10001000", "11111111", "11111111", --528
				"00000001", "00000010", "01001000", "00010000", --532
				"00100000", "10001001", "00000000", "00000000", --536
				"00100100", "10000111", "11111111", "11111011", --540
				"00000100", "00000001", "00000000", "00000000", --544
				"00000100", "00000010", "00000000", "00000000", --548
				"00000100", "00000100", "00000000", "00000000", --552
				"00000100", "00000101", "00000000", "00000000", --556
				"00000100", "00000110", "00000000", "00000011", --560
				"00000100", "00000111", "00000000", "00011010", --564
				"00000100", "00000011", "00000000", "00000000", --568
				"00000000", "00100010", "01000000", "00010000", --572
				"00011100", "01101001", "00000000", "00010100", --576
				"00000001", "00001001", "01010000", "00010000", --580
				"00010101", "01001011", "00000000", "00000011", --584
				"00011001", "01001100", "00000000", "00011101", --588
				"00000001", "01101100", "00001000", "00010011", --592
				"00100000", "01100001", "00000000", "00010100", --596
				"00000000", "00100010", "01000000", "00010000", --600
				"00011100", "10001001", "00000000", "00001010", --604
				"00000001", "00001001", "01010000", "00010000", --608
				"00000101", "01001101", "00000000", "00000000", --612
				"00001101", "00001000", "00000000", "00011111", --616
				"00000100", "00001011", "00000000", "00100000", --620
				"00000001", "01101000", "01011000", "00010001", --624
				"00000100", "00001100", "00000000", "00000000", --628
				"00101001", "10001000", "00000000", "00000011", --632
				"00010101", "01001010", "00000000", "00000001", --636
				"00000101", "10001100", "00000000", "00000001", --640
				"00110000", "00000000", "00000000", "10011110", --644
				"00000100", "00001100", "00000000", "00000000", --648
				"00101001", "10001011", "00000000", "00000011", --652
				"00011001", "10101101", "00000000", "00000001", --656
				"00000101", "10001100", "00000000", "00000001", --660
				"00110000", "00000000", "00000000", "10100011", --664
				"00000001", "01001101", "00010000", "00010011", --668
				"00100000", "10000010", "00000000", "00001010", --672
				"00000100", "10000100", "00000000", "00000001", --676
				"00001100", "10000100", "00000000", "00000011", --680
				"00000100", "01100011", "00000000", "00000001", --684
				"00100100", "01100111", "11111111", "11100010", --688
				"00000100", "10100101", "00000000", "00000001", --692
				"00100100", "10100110", "11111111", "11011110", --696
				"11111100", "00000000", "00000000", "00000000", --700 Halt 
			
				"11111100", "00000000", "00000000", "00000000", -- Halt
				"11111100", "00000000", "00000000", "00000000",-- halt repeat
				
--				"00000000", "00000000", "00000000", "00000000",	--704
--				"00000000", "00000000", "00000000", "00000000",--708
				"00000000", "00000000", "00000000", "00000000",--712
				
				"00000000", "00000000", "00000000", "00000000",--716
				"00000000", "00000000", "00000000", "00000000",--720
				"00000000", "00000000", "00000000", "00000000",--724
				"00000000", "00000000", "00000000", "00000000",--728
				"00000000", "00000000", "00000000", "00000000",--732
				"00000000", "00000000", "00000000", "00000000",--736
				"00000000", "00000000", "00000000", "00000000",--740 -- 10
				
				"00000000", "00000000", "00000000", "00000000",--744
				"00000000", "00000000", "00000000", "00000000",--748
				"00000000", "00000000", "00000000", "00000000",--752
				"00000000", "00000000", "00000000", "00000000",--760
				"00000000", "00000000", "00000000", "00000000",--764
				"00000000", "00000000", "00000000", "00000000",--768
				"00000000", "00000000", "00000000", "00000000",--772
				"00000000", "00000000", "00000000", "00000000",--776
				"00000000", "00000000", "00000000", "00000000",--780
				"00000000", "00000000", "00000000", "00000000",--784 -- 20
				
				"00000000", "00000000", "00000000", "00000000",--788
				"00000000", "00000000", "00000000", "00000000",--792
				"00000000", "00000000", "00000000", "00000000",--796
				"00000000", "00000000", "00000000", "00000000",--800
															
															
															-- Enc Begins
				"00011100", "00000001", "00000000", "00101110",--800 
				"00011100", "00000010", "00000000", "00101111",--804 
				"00011100", "00010001", "00000000", "00010100", --808
				"00011100", "00010010", "00000000", "00010101", --812
				"00000000", "00110001", "00001000", "00010000", --816
				"00000000", "01010010", "00010000", "00010000", --820
				"00000100", "00000011", "00000000", "00000001", --824
				"00000100", "00010000", "00000000", "00001101", --828
				"00000000", "00100001", "00100000", "00010100", --832
				"00000000", "01000010", "00101000", "00010100", --836
				"00000000", "00100010", "00110000", "00010100", --840
				"00000000", "10000101", "00111000", "00010100", --844
				"00000000", "11000111", "01000000", "00010100", --848
				"00000000", "00001000", "01001000", "00010000", --852
				"00001100", "01001010", "00000000", "00011111", --856
				"00000100", "00001011", "00000000", "00100000", --860
				"00000001", "01101010", "01011000", "00010001", --864
				"00000100", "00001100", "00000000", "00000000", --868
				"00101001", "10001010", "00000000", "00000011", --872
				"00010101", "00001000", "00000000", "00000001", --876
				"00000101", "10001100", "00000000", "00000001", --880
				"00110000", "00000000", "00000000", "11011010", --884
				"00000100", "00001100", "00000000", "00000000", --888
				"00101001", "10001011", "00000000", "00000011", --892
				"00011001", "00101001", "00000000", "00000001", --896
				"00000101", "10001100", "00000000", "00000001", --900
				"00110000", "00000000", "00000000", "11011111", 
				"00000001", "00001001", "01101000", "00010011", 
				"00000000", "01100011", "01110000", "00010000", 
				"00011101", "11001111", "00000000", "00010100", 
				"00000001", "10101111", "00001000", "00010000", 
				"00000000", "00100001", "00100000", "00010100", 
				"00000000", "01000010", "00101000", "00010100", 
				"00000000", "01000001", "00110000", "00010100", 
				"00000000", "10100100", "00111000", "00010100", 
				"00000000", "11100110", "01000000", "00010100", 
				"00000000", "00001000", "01001000", "00010000", 
				"00001100", "00101010", "00000000", "00011111", 
				"00000100", "00001011", "00000000", "00100000", 
				"00000001", "01101010", "01011000", "00010001", 
				"00000100", "00001100", "00000000", "00000000", 
				"00101001", "10001010", "00000000", "00000011", 
				"00010101", "00001000", "00000000", "00000001", 
				"00000101", "10001100", "00000000", "00000001", 
				"00110000", "00000000", "00000000", "11110001", 
				"00000100", "00001100", "00000000", "00000000", 
				"00101001", "10001011", "00000000", "00000011", 
				"00011001", "00101001", "00000000", "00000001", 
				"00000101", "10001100", "00000000", "00000001", 
				"00110000", "00000000", "00000000", "11110110", 
				"00000001", "00001001", "01101000", "00010011", 
				"00000000", "01100011", "01110000", "00010000", 
				"00011101", "11001111", "00000000", "00010101", 
				"00000001", "10101111", "00010000", "00010000", 
				"00000100", "01100011", "00000000", "00000001", 
				"00100100", "01110000", "11111111", "11010000",--blt 
				"00100000", "00000001", "00000000", "00110000", 
				"00100000", "00000010", "00000000", "00110001", 
				"00011100", "00010100", "00000000", "00110000", 
				"00011100", "00010101", "00000000", "00110001",
				"11111100", "00000000", "00000000", "00000000", -- Halt, addr = 1040
				"11111100", "00000000", "00000000", "00000000",-- halt repeat
				
				
				--"00000000", "00000000", "00000000", "00000000",--1040
    			--"00000000", "00000000", "00000000", "00000000",--1044

				"00000000", "00000000", "00000000", "00000000", --1048
				"00000000", "00000000", "00000000", "00000000", --1052
				"00000000", "00000000", "00000000", "00000000", --1056
				"00000000", "00000000", "00000000", "00000000", --1060
				"00000000", "00000000", "00000000", "00000000", --1064
				"00000000", "00000000", "00000000", "00000000", --1068
				"00000000", "00000000", "00000000", "00000000", --1072
				"00000000", "00000000", "00000000", "00000000", --1076
				"00000000", "00000000", "00000000", "00000000", --1080
				"00000000", "00000000", "00000000", "00000000", -- 1084/10
				
				"00000000", "00000000", "00000000", "00000000", --1088
				"00000000", "00000000", "00000000", "00000000", --1092
				"00000000", "00000000", "00000000", "00000000", --1096
				--"00000000", "00000000", "00000000", "00000000", --1100 --16
				
																				-- Dec Begins
				"00011100", "00000001", "00000000", "00110000", --1100
				"00011100", "00000010", "00000000", "00110001", --1104
				"00000100", "00000011", "00000000", "00001100", --1108
				"00000000", "01100011", "01110000", "00010000", --1112
				"00011101", "11001111", "00000000", "00010101", --1116
				"00000000", "01001111", "01000000", "00010001", --1120
				"00000000", "00001000", "01001000", "00010000", --1124
				"00001100", "00101010", "00000000", "00011111", --1128
				"00000100", "00001011", "00000000", "00100000", --1132
				"00000001", "01101010", "01011000", "00010001", --1136
				"00000100", "00001100", "00000000", "00000000", --1140
				"00101001", "10001010", "00000000", "00000011", --1144 beq
				"00011001", "00001000", "00000000", "00000001", --1148 
				"00000101", "10001100", "00000000", "00000001", --1152
				"00110000", "00000000", "00000001", "00011110", --1156
				"00000100", "00001100", "00000000", "00000000", --1160
				"00101001", "10001011", "00000000", "00000011", --1164 beq
				"00010101", "00101001", "00000000", "00000001", --1168
				"00000101", "10001100", "00000000", "00000001", --1172
				"00110000", "00000000", "00000001", "00100011", --1176
				"00000001", "00001001", "01101000", "00010011", --1180
				"00000000", "00100001", "00100000", "00010100", --1184
				"00000001", "10101101", "00101000", "00010100", --1188
				"00000001", "10100001", "00110000", "00010100", --1192
				"00000000", "10100100", "00111000", "00010100", --1196
				"00000000", "11100110", "00010000", "00010100", --1200
				"00000000", "01100011", "01110000", "00010000", --1204
				"00011101", "11001111", "00000000", "00010100", --1208
				"00000000", "00101111", "01000000", "00010001", --1212
				"00000000", "00001000", "01001000", "00010000", --1216
				"00001100", "01001010", "00000000", "00011111", --1220
				"00000100", "00001011", "00000000", "00100000", --1224
				"00000001", "01101010", "01011000", "00010001", --1228
				"00000100", "00001100", "00000000", "00000000", --1232
				"00101001", "10001010", "00000000", "00000011", --1236--beq
				"00011001", "00001000", "00000000", "00000001", --1240
				"00000101", "10001100", "00000000", "00000001", --1244
				"00110000", "00000000", "00000001", "00110101", --1248
				"00000100", "00001100", "00000000", "00000000", --1252
				"00101001", "10001011", "00000000", "00000011", --1256--beq
				"00010101", "00101001", "00000000", "00000001", --1260
				"00000101", "10001100", "00000000", "00000001", --1264
				"00110000", "00000000", "00000001", "00111010", --1268
				"00000001", "00001001", "01101000", "00010011", --1272
				"00000001", "10101101", "00100000", "00010100", --1276
				"00000000", "01000010", "00101000", "00010100", --1280
				"00000001", "10100010", "00110000", "00010100", --1284
				"00000000", "10000101", "00111000", "00010100", --1288
				"00000000", "11000111", "00001000", "00010100", --1292
				"00001000", "01100011", "00000000", "00000001", --1296
				"00101100", "01100000", "11111111", "11010000", --1300--bne
				"00011100", "00010001", "00000000", "00010100", 
				"00011100", "00010010", "00000000", "00010101", 
				"00000000", "00110001", "00001000", "00010001", 
				"00000000", "01010010", "00010000", "00010001", 
				"00100000", "00000001", "00000000", "00110000", 
				"00100000", "00000010", "00000000", "00110001", 
				"11111100", "00000000", "00000000", "00000000", -- Halt, addr = 1328
				"11111100", "00000000", "00000000", "00000000", -- 1332
				"00000000", "00000000", "00000000", "00000000"); -- 1336

  
				
--				"00000100", "00000001", "00000000", "00000111", --ADDI R1, R0, 7 // R1 = 7
--				"00000100", "00000010", "00000000", "00001000", --ADDI R2, R0, 8 // R2 = 8
--				"00000000", "01000001", "00011000", "00010000", --ADD R3, R1, R2 // R3 = R1 + R2 =15
--				"11111100", "00000000", "00000000", "00000000"); -- Halt
				
				
				
--			
--				
--				"00110000", "00000000", "00000001", "00000100",		--location 0
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				"00000000", "00000000", "00000000", "00000000",
--				--store p and q
--				"00000100", "00000001", "10110111", "11100001",	--	ADDI R0 R1 0xB7E1  location 460
--				"00010100", "00100010", "00000000", "00010000",	--SHL R1 R2 0x0010
--				"00000100", "00000011", "01010001", "01100011",	--ADDI R0 R3 0x5163
--				"00000000", "01000011", "00100000", "00010011",	--OR R2 R3 R4
--				"00100000", "00000100", "00000000", "00001110",	--SW R0 R4 0x000E
--				"00000100", "00000101", "10011110", "00110111",	--ADDI R0 R5 0x9E37
--				"00010100", "10100110", "00000000", "00010000",	-- SHL R5 R6 0x0010
--				"00000100", "00000111", "01111001", "10111001",	--ADDI R0 R7 0x79B9
--				"00000000", "11000111", "01000000", "00010011",	--OR R6 R7 R8
--				"00100000", "00001000", "00000000", "00001111",		--SW R0 R8 0x000F--location 496
--				
----key gen		
--"00011100","00000001","00000000","00001110",	--Lw R0, R1, 14		// R1 = P
--"00011100","00000010","00000000","00001111",	--Lw R0, R2, 15		// R2 = Q
--"00000100","00000100","00000000","00010100",	--Addi R0, R4, 20		// R4 = 20
--"00100000","10000001","00000000","00000000",	--Sw R4, R1, 0		// S[0] = P
--"00000100","00000110","00000000","00011001",	--Addi R0, R6, 25		// Initializing R6 = 25
--"00000000","10000110","00111000","00010000",	--Add R4, R6, R7		// R7 = 46 // End  
--"00000100","10000100","00000000","00000001",	--Addi R4, R4, 1		// increment i
--"00011100","10001000","11111111","11111111",	--Lw R4, R8, 0xFFFF	// S[ i - 1 ] 	
--"00000001","00000010","01001000","00010000",	--add R8, R2, R9		// R9 = R2 + R8 
--"00100000","10001001","00000000","00000000",	-- Sw R4, R9, 0		// S[i] = S[i-1] + Q 
--"00100100","10000111","00000010","00001100",	--BLT R4, R7, LoopKeyInit	 
--"00000100","00000001","00000000","00000000",	--Addi R0, R1, 0		// Initialize A = 0
--"00000100","00000010","00000000","00000000",	--Addi R0, R2, 0		// Initialize B = 0
--"00000100","00000100","00000000","00000000",	--Addi R0, R4, 0		// Initialize j = 0
--"00000100","00000101","00000000","00000000",	--Addi R0, R5, 0 		// Initialize k = 0
--"00000100","00000110","00000000","00000011",	--Addi R0, R6, 3 		// Outer loop count
--"00000100","00000111","00000000","00011010",	--Addi R0, R7, 26		// Inner loop count
--"00000100","00000011","00000000","00000000",	--Addi R0, R3, 0		//Initialize i = 0
--"00000000","00100010","01000000","00010000",	--Add R1, R2, R8		// A+B
--"00011100","01101001","00000000","00010100",	--Lw R3, R9, 20		// S[i]
--"00000000","01001001","01010000","00010000",	--Add R2, R9, R10		// S[i] + (A+B)
--"00010101","01001011","00000000","00000011",	--SHL R10, R11, 3		// R11 = R10 << 3
--"00011001","01001100","00000000","00011101",	--SHR R10, R12, 29	// R12 = R10 >> 29
--"00000001","01101100","00001000","00010011",	--OR R11, R12, R1		// A = R11 OR R12 
--"00100000","01100001","00000000","00010100",	--Sw R3, R1, 20		// S[i] = A
--"00000000","00100010","01000000","00010000",	--Add R1, R2, R8		// A+B
--"00011100","10001001","00000000","00001010", --Lw R4, R9, 10		// L[j]
--"00000001","00001001","01010000","00010000",	--Add R8, R9, R10		// L[j] + (A+B)
--"00000101","01001101","00000000","00000000",	--Addi R10, R13, 0	// copy of R10	
--"00001101","00001000","00000000","00011111",	--ANDI R8, R8, 0x0000001F//mod 32 of (A+B)//Left Shift --Amount
--"00000100","00001011","00000000","00100000",	--Addi R0, R11, 32	
--"00000001","01101000","01011000","00010000",	--Sub R11, R8, R11// R11= 32-R8		// Right --Shift Amount
--			--// Data Dependent Circular Left Rotate begins
--"00000100","00001100","00000000","00000000",	--Addi R0, R12, 0		// Initializing R12  
----LoopSHL: 
--"00101001","10001000","00000010","10001000",	--BEQ R12, R8, EndLoopSHL  
--"00010101","01001010","00000000","00000001",	--SHL R10, R10, 1		
--"00000101","10001100","00000000","00000001",	--Addi R12, R12, 1	// Incrementing R12
--"00110000","00000000","00000010","01111000",		--Jmp LoopSHL
----EndLoopSHL:
--"00000100","00001100","00000000","00000000",	--Addi R0, R12, 0		// Initializing R12  
----LoopSHR: 
--"00101001","10001011","00000010","10011100",	--BEQ R12, R11, EndLoopSHR  
--"00011001","10101101","00000000","00000001",	--SHR R13, R13, 1	
--"00000101","10001100","00000000","00000001",	--Addi R12, R12, 1	// Incrementing R12
--"00110000","00000000","00000010","10001100",	--Jmp LoopSHR
----EndLoopSHR:
--"00000001","01001101","00010000","00010011",	--OR R10, R13, R2	// B = R10 OR R13// Result of -----Data Dependent Circular Left Rotate
--"00100000","10000010","00000000","00001010",	--Sw R4, R2, 10		// L[j] = B	
--"00000100","10000100","00000000","00000001",	--Addi R4, R4, 1		//Increment j
--"00000100","10000100","00000000","00000011",	--ANDI R4, R4, 0x00000003	//Mod 4 of j
--"00000100","01100011","00000000","00000001",	--Addi R3, R3,1		// Increment i
--"00100100","01100111","00000010","00111100",	 --BLT R3, R7, LoopKeyExp2
--"00000100","10100101","00000000","00000001",	--Addi R5, R5, 1		// Increment k
--"00100100","10100110","00000010","00111000",	--BLT R5, R6, LoopKeyExp1
--"11111100","00000000","00000000","00000000"


--"00000100", "00000001", "00000000", "00000010", --ADDI R1, R0, 2 //R1=R0+2(decimal)
--				"00000100", "00000011", "00000000", "00001010", --ADDI R3, R0, 10 //R3=R0+10(decimal)
--				"00000100", "00000100", "00000000", "00001110", --ADDI R4, R0, 14 //R4=R0+14(decimal)
--				"00000100", "00000101", "00000000", "00000010", --ADDI R5, R0, 2 //R5=R0+2
--				"00100000", "01100100", "00000000", "00000010", --SW R4, 2(R3) //Mem[R3+2]=R4
--				"00100000", "01100011", "00000000", "00000001", --SW R3, 1(R3) //Mem[R3+1]=R3
--				"00000000", "10000011", "00100000", "00010001", --SUB R4, R4, R3 //R4=R4-R3
--				"00001000", "00000100", "00000000", "00000001", --SUBI R4, R0, 1 //R4=R0-1(decimal)
--				"00000000", "01100010", "00100000", "00010010", --AND R4, R2, R3 //R4=R2 and R3
--				"00001100", "01000100", "00000000", "00001010", --ANDI R4, R2, 10 //R4=R2 and 10(decimal)
--				"00000000", "01100010", "00100000", "00010011", --OR R4, R2, R3 //R4= R2 or R3
--				"00011100", "01100010", "00000000", "00000001", --LW R2, 1(R3) //R2=Mem[1+R3]
--				"00010000", "01000100", "00000000", "00001010", --ORI R4, R2, 10 //R4=R2 or 10(decimal)
--				"00000000", "01100010", "00100000", "00010100", --NOR R4, R2, R3 //R4= R2 nor R3
--				"00010100", "01000100", "00000000", "00001010", --SHL R4, R2, 10 //R4= R2 << 10(decimal)
--				"00011000", "01000100", "00000000", "00001010", --SHR R4, R2, 10 //R4=R2 >> 10(decimal)
--				"00101000", "00000101", "11111111", "11111110", --BEQ R5, R0, -2
--				"00100100", "10000101", "00000000", "00000000", --BLT R5, R4, 0
--				"00101100", "10000101", "00000000", "00000000", --BNE R5, R4, 0
--				"00110000", "00000000", "00000000", "00010100", --JMP 20
--				"11111100", "00000000", "00000000", "00000000"); --HAL
   

BEGIN
 -- imem[PC] & imem[PC+1] & imem[PC+2] & imem[PC+3]
  Instruction<=imem(CONV_INTEGER(PC)) & imem(CONV_INTEGER(PC)+1) & 
					imem(CONV_INTEGER(PC)+2) & imem(CONV_INTEGER(PC)+3);
END rtl;